//behavioral model.
//8 bit adder using full adder more specifically, this is a ripple carry adder.

//import full adder file, which is already created.
`include "fullAdder.v"

//starting module.
module ebaUfa(a,b,cin,sum,cout);

// i/o declaration.
input [7:0]a;
input [7:0]b;
input cin;
output [7:0]sum;
output cout;

// intermediate value declaration.
wire [6:0]c;

//Full adder one.
fullAdder a1(a[0],b[0],cin,sum[0],c[0]);
//Full adder two.
fullAdder a2(a[1],b[1],c[0],sum[1],c[1]);
//Full adder three.
fullAdder a3(a[2],b[2],c[1],sum[2],c[2]);
//Full adder four.
fullAdder a4(a[3],b[3],c[2],sum[3],c[3]);
//Full adder five.
fullAdder a5(a[4],b[4],c[3],sum[4],c[4]);
//Full adder six.
fullAdder a6(a[5],b[5],c[4],sum[5],c[5]);
//Full adder seven.
fullAdder a7(a[6],b[6],c[5],sum[6],c[6]);
//Full adder eight.
fullAdder a8(a[7],b[7],c[6],sum[7],cout);

//module finished.
endmodule
